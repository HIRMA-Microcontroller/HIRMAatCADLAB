library verilog;
use verilog.vl_types.all;
entity aftab_testbench is
end aftab_testbench;
