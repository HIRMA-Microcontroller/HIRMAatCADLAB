library verilog;
use verilog.vl_types.all;
entity aftab_AAU_TB is
end aftab_AAU_TB;
