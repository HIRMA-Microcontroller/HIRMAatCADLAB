library verilog;
use verilog.vl_types.all;
entity aftab_sgn_divider_TB is
end aftab_sgn_divider_TB;
