library verilog;
use verilog.vl_types.all;
entity aftab_DAWU_TB is
end aftab_DAWU_TB;
