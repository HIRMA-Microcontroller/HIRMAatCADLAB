library verilog;
use verilog.vl_types.all;
entity collection_tb is
end collection_tb;
