library verilog;
use verilog.vl_types.all;
entity aftab_boothTB is
end aftab_boothTB;
