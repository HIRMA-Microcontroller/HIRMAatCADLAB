library verilog;
use verilog.vl_types.all;
entity MCU_TB is
end MCU_TB;
