library verilog;
use verilog.vl_types.all;
entity aftab_divider_TB is
end aftab_divider_TB;
