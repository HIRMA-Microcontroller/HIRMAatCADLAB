library verilog;
use verilog.vl_types.all;
entity aftab_datapath is
    generic(
        size            : integer := 32
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        writeRegFile    : in     vl_logic;
        setOne          : in     vl_logic;
        setZero         : in     vl_logic;
        compareSignedUnsignedBar: in     vl_logic;
        selPC           : in     vl_logic;
        selI4           : in     vl_logic;
        selAdd          : in     vl_logic;
        selJL           : in     vl_logic;
        selADR          : in     vl_logic;
        selPCJ          : in     vl_logic;
        selInc4PC       : in     vl_logic;
        selBSU          : in     vl_logic;
        selLLU          : in     vl_logic;
        selASU          : in     vl_logic;
        selAAU          : in     vl_logic;
        selDARU         : in     vl_logic;
        selP1           : in     vl_logic;
        selP2           : in     vl_logic;
        selImm          : in     vl_logic;
        ldPC            : in     vl_logic;
        zeroPC          : in     vl_logic;
        ldADR           : in     vl_logic;
        zeroADR         : in     vl_logic;
        ldDR            : in     vl_logic;
        zeroDR          : in     vl_logic;
        ldIR            : in     vl_logic;
        zeroIR          : in     vl_logic;
        ldByteSigned    : in     vl_logic;
        ldHalfSigned    : in     vl_logic;
        load            : in     vl_logic;
        selShift        : in     vl_logic_vector(1 downto 0);
        addSubBar       : in     vl_logic;
        pass            : in     vl_logic;
        selAuipc        : in     vl_logic;
        muxCode         : in     vl_logic_vector(11 downto 0);
        selLogic        : in     vl_logic_vector(1 downto 0);
        startDAWU       : in     vl_logic;
        startDARU       : in     vl_logic;
        startMultiplyAAU: in     vl_logic;
        startDivideAAU  : in     vl_logic;
        signedSigned    : in     vl_logic;
        signedUnsigned  : in     vl_logic;
        unsignedUnsigned: in     vl_logic;
        selAAL          : in     vl_logic;
        selAAH          : in     vl_logic;
        dataInstrBar    : in     vl_logic;
        nBytes          : in     vl_logic_vector(1 downto 0);
        memReady        : in     vl_logic;
        memDataIn       : in     vl_logic_vector(7 downto 0);
        memDataOut      : out    vl_logic_vector(7 downto 0);
        memAddrDAWU     : out    vl_logic_vector;
        memAddrDARU     : out    vl_logic_vector;
        writeMem        : out    vl_logic;
        readMem         : out    vl_logic;
        IR              : out    vl_logic_vector;
        lt              : out    vl_logic;
        eq              : out    vl_logic;
        gt              : out    vl_logic;
        completeDAWU    : out    vl_logic;
        completeDARU    : out    vl_logic;
        completeAAU     : out    vl_logic;
        selCSR          : in     vl_logic;
        machineExternalInterrupt: in     vl_logic;
        machineTimerInterrupt: in     vl_logic;
        machineSoftwareInterrupt: in     vl_logic;
        userExternalInterrupt: in     vl_logic;
        userTimerInterrupt: in     vl_logic;
        userSoftwareInterrupt: in     vl_logic;
        platformInterruptSignals: in     vl_logic_vector(15 downto 0);
        ldValueCSR      : in     vl_logic_vector(2 downto 0);
        mipCCLdDisable  : in     vl_logic;
        selImmCSR       : in     vl_logic;
        selP1CSR        : in     vl_logic;
        selReadWriteCSR : in     vl_logic;
        clrCSR          : in     vl_logic;
        setCSR          : in     vl_logic;
        selPC_CSR       : in     vl_logic;
        selTval_CSR     : in     vl_logic;
        selMedeleg_CSR  : in     vl_logic;
        selMideleg_CSR  : in     vl_logic;
        selCCMip_CSR    : in     vl_logic;
        selCause_CSR    : in     vl_logic;
        selMepc_CSR     : in     vl_logic;
        selInterruptAddressDirect: in     vl_logic;
        selInterruptAddressVectored: in     vl_logic;
        writeRegBank    : in     vl_logic;
        dnCntCSR        : in     vl_logic;
        upCntCSR        : in     vl_logic;
        ldCntCSR        : in     vl_logic;
        zeroCntCSR      : in     vl_logic;
        ldFlags         : in     vl_logic;
        zeroFlags       : in     vl_logic;
        ldDelegation    : in     vl_logic;
        ldMachine       : in     vl_logic;
        ldUser          : in     vl_logic;
        loadMieReg      : in     vl_logic;
        loadMieUieField : in     vl_logic;
        mirrorUser      : in     vl_logic;
        machineStatusAlterationPreCSR: in     vl_logic;
        userStatusAlterationPreCSR: in     vl_logic;
        machineStatusAlterationPostCSR: in     vl_logic;
        userStatusAlterationPostCSR: in     vl_logic;
        checkMisalignedDARU: in     vl_logic;
        checkMisalignedDAWU: in     vl_logic;
        selCSRAddrFromInst: in     vl_logic;
        selRomAddress   : in     vl_logic;
        ecallFlag       : in     vl_logic;
        illegalInstrFlag: in     vl_logic;
        instrMisalignedOut: out    vl_logic;
        loadMisalignedOut: out    vl_logic;
        storeMisalignedOut: out    vl_logic;
        dividedByZeroOut: out    vl_logic;
        validAccessCSR  : out    vl_logic;
        readOnlyCSR     : out    vl_logic;
        mirror          : out    vl_logic;
        ldMieReg        : out    vl_logic;
        ldMieUieField   : out    vl_logic;
        interruptRaise  : out    vl_logic;
        exceptionRaise  : out    vl_logic;
        delegationMode  : out    vl_logic_vector(1 downto 0);
        previousPRV     : out    vl_logic_vector(1 downto 0);
        modeTvec        : out    vl_logic_vector(1 downto 0)
    );
end aftab_datapath;
