`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/28/2023 09:54:51 AM
// Design Name: 
// Module Name: auto_fifo_fill
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module auto_fifo_fill
#(parameter fifo_depth = 2000)
(
	input clk,
	input rst,
	input start,
	output reg direct_fifo,
	output reg [7:0] direct_buf_in,
	output reg direct_wr_en_buf
    );
	
	parameter BUF_SIZE = fifo_depth;
	integer i;
	
	reg [7:0] mem [0: BUF_SIZE-1];
	
	reg [3:0] ps, ns;
	
	reg [31:0] cnt;
	reg cen;
	reg init0;
	
	localparam [3:0] IDLE = 0,
					         INIT = 1,
					         PASS = 2,
					         END  = 3;
	
	always @(posedge clk) begin
	
		if(rst) begin
			for(i=0; i<BUF_SIZE; i=i+1) begin
				mem[i] <= 0;
			end
			mem[0 ] <=	8'b00001111;
			mem[1 ] <=	8'b10110011;
			mem[2 ] <=	8'b00000000;
			mem[3 ] <=	8'b00000000;
			mem[4 ] <=	8'b00000000;
			mem[5 ] <=	8'b00010011;
			mem[6 ] <=	8'b00000001;
			mem[7 ] <=	8'b00010000;
			mem[8 ] <=	8'b00000000;
			mem[9 ] <=	8'b10010011;
			mem[10] <=	8'b00000001;
			mem[11] <=	8'b01010000;
			mem[12] <=	8'b00000000;
			mem[13] <=	8'b00010011;
			mem[14] <=	8'b00000010;
			mem[15] <=	8'b00010000;
			mem[16] <=	8'b00000000;
			mem[17] <=	8'b01100011;
			mem[18] <=	8'b10001010;
			mem[19] <=	8'b00110000;
			mem[20] <=	8'b00000000;
			mem[21] <=	8'b00110011;
			mem[22] <=	8'b00000010;
			mem[23] <=	8'b01000001;
			mem[24] <=	8'b00000010;
			mem[25] <=	8'b00010011;
			mem[26] <=	8'b00000001;
			mem[27] <=	8'b00010001;
			mem[28] <=	8'b00000000;
			mem[29] <=	8'b10010011;
			mem[30] <=	8'b10000000;
			mem[31] <=	8'b00010000;
			mem[32] <=	8'b00000000;
			mem[33] <=	8'b11101111;
			mem[34] <=	8'b11110010;
			mem[35] <=	8'b00011111;
			mem[36] <=	8'b11111111;
			mem[37] <=	8'b00010011;
			mem[38] <=	8'b00000011;
			mem[39] <=	8'b00100000;
			mem[40] <=	8'b00000001;
			mem[41] <=	8'b10110011;
			mem[42] <=	8'b01000011;
			mem[43] <=	8'b01100010;
			mem[44] <=	8'b00000010;
			mem[45] <=	8'b00110011;
			mem[46] <=	8'b01100100;
			mem[47] <=	8'b01100010;
			mem[48] <=	8'b00000010;
			mem[49] <=	8'b00100011;
			mem[50] <=	8'b00100000;
			mem[51] <=	8'b01110000;
			mem[52] <=	8'b00100000;
			mem[53] <=	8'b00010011;
			mem[54] <=	8'b00001010;
			mem[55] <=	8'b00000000;
			mem[56] <=	8'b01000000;
			mem[57] <=	8'b00010011;
			mem[58] <=	8'b00011010;
			mem[59] <=	8'b00101010;
			mem[60] <=	8'b00000000;
			mem[61] <=	8'b00100011;
			mem[62] <=	8'b00100000;
			mem[63] <=	8'b01111010;
			mem[64] <=	8'b00000000;
			mem[65] <=	8'b00000011;
			mem[66] <=	8'b00100101;
			mem[67] <=	8'b00001010;
			mem[68] <=	8'b00000000;
			mem[69] <=	8'b00010011;
			mem[70] <=	8'b00011010;
			mem[71] <=	8'b00001010;
			mem[72] <=	8'b00000001;
			mem[73] <=	8'b10110011;
			mem[74] <=	8'b00001010;
			mem[75] <=	8'b00001010;
			mem[76] <=	8'b00000000;
			mem[77] <=	8'b00010011;
			mem[78] <=	8'b01011010;
			mem[79] <=	8'b00011010;
			mem[80] <=	8'b00000000;
			mem[81] <=	8'b10110011;
			mem[82] <=	8'b00001010;
			mem[83] <=	8'b01011010;
			mem[84] <=	8'b00000001;
			mem[85] <=	8'b00010011;
			mem[86] <=	8'b01011010;
			mem[87] <=	8'b00101010;
			mem[88] <=	8'b00000000;
			mem[89] <=	8'b10110011;
			mem[90] <=	8'b00001010;
			mem[91] <=	8'b01011010;
			mem[92] <=	8'b00000001;
			mem[93] <=	8'b00010011;
			mem[94] <=	8'b01011010;
			mem[95] <=	8'b01011010;
			mem[96] <=	8'b00000000;
			mem[97] <=	8'b10110011;
			mem[98] <=	8'b00001010;
			mem[99] <=	8'b01011010;
			mem[100] <=	8'b00000001;
			mem[101] <=	8'b00010011;
			mem[102] <=	8'b01011010;
			mem[103] <=	8'b01011010;
			mem[104] <=	8'b00000000;
			mem[105] <=	8'b10110011;
			mem[106] <=	8'b00001010;
			mem[107] <=	8'b01011010;
			mem[108] <=	8'b00000001;
			mem[109] <=	8'b00010011;
			mem[110] <=	8'b01011010;
			mem[111] <=	8'b00011010;
			mem[112] <=	8'b00000000;
			mem[113] <=	8'b10110011;
			mem[114] <=	8'b00001010;
			mem[115] <=	8'b01011010;
			mem[116] <=	8'b00000001;
			mem[117] <=	8'b00010011;
			mem[118] <=	8'b01011010;
			mem[119] <=	8'b00011010;
			mem[120] <=	8'b00000000;
			mem[121] <=	8'b10110011;
			mem[122] <=	8'b00001010;
			mem[123] <=	8'b01011010;
			mem[124] <=	8'b00000001;
			mem[125] <=	8'b00010011;
			mem[126] <=	8'b00001011;
			mem[127] <=	8'b11110000;
			mem[128] <=	8'b01111111;
			mem[129] <=	8'b00010011;
			mem[130] <=	8'b00011011;
			mem[131] <=	8'b00101011;
			mem[132] <=	8'b00000000;
			mem[133] <=	8'b10110011;
			mem[134] <=	8'b00001010;
			mem[135] <=	8'b01011011;
			mem[136] <=	8'b00000001;
			mem[137] <=	8'b10010011;
			mem[138] <=	8'b10001010;
			mem[139] <=	8'b11001010;
			mem[140] <=	8'b11111110;
			mem[141] <=	8'b10010011;
			mem[142] <=	8'b00001001;
			mem[143] <=	8'b11110000;
			mem[144] <=	8'b00001111;
			mem[145] <=	8'b00100011;
			mem[146] <=	8'b10100000;
			mem[147] <=	8'b00111010;
			mem[148] <=	8'b00000001;
			mem[149] <=	8'b10010011;
			mem[150] <=	8'b10001010;
			mem[151] <=	8'b01001010;
			mem[152] <=	8'b00000000;
			mem[153] <=	8'b10010011;
			mem[154] <=	8'b00001001;
			mem[155] <=	8'b11110000;
			mem[156] <=	8'b00011111;
			mem[157] <=	8'b00100011;
			mem[158] <=	8'b10100000;
			mem[159] <=	8'b00111010;
			mem[160] <=	8'b00000001;
			mem[161] <=	8'b10010011;
			mem[162] <=	8'b10001010;
			mem[163] <=	8'b01001010;
			mem[164] <=	8'b00000000;
			mem[165] <=	8'b10010011;
			mem[166] <=	8'b00001001;
			mem[167] <=	8'b00100000;
			mem[168] <=	8'b00000000;
			mem[169] <=	8'b00100011;
			mem[170] <=	8'b10000000;
			mem[171] <=	8'b00111010;
			mem[172] <=	8'b00000001;
			mem[173] <=	8'b10010011;
			mem[174] <=	8'b00001001;
			mem[175] <=	8'b01010000;
			mem[176] <=	8'b00000000;
			mem[177] <=	8'b00100011;
			mem[178] <=	8'b10000000;
			mem[179] <=	8'b00111010;
			mem[180] <=	8'b00000001;
			mem[181] <=	8'b00000011;
			mem[182] <=	8'b10001001;
			mem[183] <=	8'b00001010;
			mem[184] <=	8'b00000000;
			mem[185] <=	8'b10010011;
			mem[186] <=	8'b10001010;
			mem[187] <=	8'b10001010;
			mem[188] <=	8'b11111110;
			mem[189] <=	8'b10010011;
			mem[190] <=	8'b00001011;
			mem[191] <=	8'b00100000;
			mem[192] <=	8'b00011011;
			mem[193] <=	8'b00100011;
			mem[194] <=	8'b10100000;
			mem[195] <=	8'b01111010;
			mem[196] <=	8'b00000001;
			mem[197] <=	8'b10010011;
			mem[198] <=	8'b10001010;
			mem[199] <=	8'b10001010;
			mem[200] <=	8'b00000000;
			mem[201] <=	8'b00010011;
			mem[202] <=	8'b00001100;
			mem[203] <=	8'b10010000;
			mem[204] <=	8'b00001010;
			mem[205] <=	8'b00100011;
			mem[206] <=	8'b10000000;
			mem[207] <=	8'b10001010;
			mem[208] <=	8'b00000001;
			mem[209] <=	8'b00010011;
			mem[210] <=	8'b00001100;
			mem[211] <=	8'b00010000;
			mem[212] <=	8'b00000000;
			mem[213] <=	8'b10010011;
			mem[214] <=	8'b10001010;
			mem[215] <=	8'b01001010;
			mem[216] <=	8'b00000000;
			mem[217] <=	8'b00100011;
			mem[218] <=	8'b10000000;
			mem[219] <=	8'b10001010;
			mem[220] <=	8'b00000001;
			mem[221] <=	8'b00010011;
			mem[222] <=	8'b00001100;
			mem[223] <=	8'b11100000;
			mem[224] <=	8'b00000001;
			mem[225] <=	8'b00100011;
			mem[226] <=	8'b10000000;
			mem[227] <=	8'b10001010;
			mem[228] <=	8'b00000001;
			mem[229] <=	8'b10010011;
			mem[230] <=	8'b10001010;
			mem[231] <=	8'b10001010;
			mem[232] <=	8'b11111111;
			mem[233] <=	8'b10000011;
			mem[234] <=	8'b10001000;
			mem[235] <=	8'b00001010;
			mem[236] <=	8'b00000000;
			
			mem[255] <=	8'b01110001;
			mem[256] <=	8'b01001001;
			
			mem[511] <=	8'h0A;
			mem[512] <=	8'h0B;
			
			mem[767] <=	8'h0C;
			mem[768] <=	8'h0D;
			
			mem[1023] <=	8'h0E;
			mem[1024] <=	8'h0F;
			
			mem[1279] <=	8'h0A;
			mem[1280] <=	8'h0B;
			
			mem[1535] <=	8'h0C;
			mem[1536] <=	8'h0D;
			
			mem[4095] <=	8'h0E;
			mem[4096] <=	8'h2F;
			
			
			mem[4999] <= 8'b10100101;
		end
		
		else begin
			for(i=0; i<BUF_SIZE; i=i+1) begin
				mem[i] <= mem[i];
			end
		end
	
	end
	
	always @(posedge clk) begin
		if(rst)
			ps <= IDLE;
			
		else
			ps <= ns;
	
	end
	
	always @(ps, start, cnt) begin
		case(ps) 
			IDLE :	ns = (start) ? INIT : IDLE;
			INIT :  ns = (!start) ? PASS : INIT;
			PASS :  ns = (cnt == BUF_SIZE) ? END : PASS;
			END  :  ns = END;
		endcase
	end
	
	always @(ps, cnt) begin
		init0 = 0;
		direct_fifo = 0;
		direct_wr_en_buf = 0;
		case(ps)
			IDLE : begin   
			end
			
			INIT : begin
				init0 = 1;
			end
			
			PASS : begin
				direct_fifo = 1;
				direct_wr_en_buf = 1;
				direct_buf_in = mem[cnt];
				cen = 1;
			end
			
			END : begin
			end
			
		endcase
		
	end
	
	
	always @(posedge clk) begin
		if(rst)
			cnt <= 0;
		else if(init0)
			cnt <= 0;
		else if(cen)
			cnt <= cnt + 1;
		else	
			cnt <= cnt;
	end
	
endmodule

