library verilog;
use verilog.vl_types.all;
entity aftab_BSU_TB is
end aftab_BSU_TB;
