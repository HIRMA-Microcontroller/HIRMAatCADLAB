library verilog;
use verilog.vl_types.all;
entity aftab_controller is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        completeDARU    : in     vl_logic;
        completeDAWU    : in     vl_logic;
        completeAAU     : in     vl_logic;
        lt              : in     vl_logic;
        eq              : in     vl_logic;
        gt              : in     vl_logic;
        IR              : in     vl_logic_vector(31 downto 0);
        interruptRaise  : in     vl_logic;
        exceptionRaise  : in     vl_logic;
        instrMisalignedOut: in     vl_logic;
        loadMisalignedOut: in     vl_logic;
        storeMisalignedOut: in     vl_logic;
        dividedByZeroOut: in     vl_logic;
        validAccessCSR  : in     vl_logic;
        readOnlyCSR     : in     vl_logic;
        mirror          : in     vl_logic;
        ldMieReg        : in     vl_logic;
        ldMieUieField   : in     vl_logic;
        delegationMode  : in     vl_logic_vector(1 downto 0);
        previousPRV     : in     vl_logic_vector(1 downto 0);
        modeTvec        : in     vl_logic_vector(1 downto 0);
        muxCode         : out    vl_logic_vector(11 downto 0);
        nBytes          : out    vl_logic_vector(1 downto 0);
        selLogic        : out    vl_logic_vector(1 downto 0);
        selShift        : out    vl_logic_vector(1 downto 0);
        selPC           : out    vl_logic;
        selI4           : out    vl_logic;
        selP1           : out    vl_logic;
        selP2           : out    vl_logic;
        selJL           : out    vl_logic;
        selADR          : out    vl_logic;
        selPCJ          : out    vl_logic;
        selImm          : out    vl_logic;
        selAdd          : out    vl_logic;
        selInc4PC       : out    vl_logic;
        selBSU          : out    vl_logic;
        selLLU          : out    vl_logic;
        selASU          : out    vl_logic;
        selAAU          : out    vl_logic;
        selDARU         : out    vl_logic;
        dataInstrBar    : out    vl_logic;
        writeRegFile    : out    vl_logic;
        addSubBar       : out    vl_logic;
        pass            : out    vl_logic;
        selAuipc        : out    vl_logic;
        comparedsignedunsignedbar: out    vl_logic;
        ldIR            : out    vl_logic;
        ldADR           : out    vl_logic;
        ldPC            : out    vl_logic;
        ldDr            : out    vl_logic;
        ldByteSigned    : out    vl_logic;
        ldHalfSigned    : out    vl_logic;
        load            : out    vl_logic;
        setOne          : out    vl_logic;
        setZero         : out    vl_logic;
        startDARU       : out    vl_logic;
        startDAWU       : out    vl_logic;
        startMultiplyAAU: out    vl_logic;
        startDivideAAU  : out    vl_logic;
        signedSigned    : out    vl_logic;
        signedUnsigned  : out    vl_logic;
        unsignedUnsigned: out    vl_logic;
        selAAL          : out    vl_logic;
        selAAH          : out    vl_logic;
        ecallFlag       : out    vl_logic;
        illegalInstrFlag: out    vl_logic;
        mipCCLdDisable  : out    vl_logic;
        selCCMip_CSR    : out    vl_logic;
        selCause_CSR    : out    vl_logic;
        selPC_CSR       : out    vl_logic;
        selTval_CSR     : out    vl_logic;
        selMedeleg_CSR  : out    vl_logic;
        selMideleg_CSR  : out    vl_logic;
        ldValueCSR      : out    vl_logic_vector(2 downto 0);
        ldCntCSR        : out    vl_logic;
        dnCntCSR        : out    vl_logic;
        upCntCSR        : out    vl_logic;
        ldFlags         : out    vl_logic;
        zeroFlags       : out    vl_logic;
        ldDelegation    : out    vl_logic;
        ldMachine       : out    vl_logic;
        ldUser          : out    vl_logic;
        loadMieReg      : out    vl_logic;
        loadMieUieField : out    vl_logic;
        mirrorUser      : out    vl_logic;
        selCSR          : out    vl_logic;
        selP1CSR        : out    vl_logic;
        selReadWriteCSR : out    vl_logic;
        selImmCSR       : out    vl_logic;
        setCSR          : out    vl_logic;
        clrCSR          : out    vl_logic;
        writeRegBank    : out    vl_logic;
        selCSRAddrFromInst: out    vl_logic;
        selRomAddress   : out    vl_logic;
        selMepc_CSR     : out    vl_logic;
        selInterruptAddressDirect: out    vl_logic;
        selInterruptAddressVectored: out    vl_logic;
        checkMisalignedDARU: out    vl_logic;
        checkMisalignedDAWU: out    vl_logic;
        machineStatusAlterationPreCSR: out    vl_logic;
        userStatusAlterationPreCSR: out    vl_logic;
        machineStatusAlterationPostCSR: out    vl_logic;
        userStatusAlterationPostCSR: out    vl_logic;
        zeroCntCSR      : out    vl_logic
    );
end aftab_controller;
