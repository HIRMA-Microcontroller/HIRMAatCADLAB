//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM, INC.
//Copyright (c) 2002-2009 ARM, Inc.
//The confidential and proprietary information contained in this file
//may only be used by a person authorised under and to the extent
//permitted by a subsisting licensing agreement from ARM Limited.
//
//(C) COPYRIGHT 2004-2009 ARM Limited.
//ALL RIGHTS RESERVED
//
//This entire notice must be reproduced on all copies of this file
//and copies of this file may only be made by a person if such person
//is permitted to do so under the terms of a subsisting license
//agreement from ARM Limited.
//

`define ARM_PROP_DELAY 1.0
`define ARM_PERIOD 1.0
`define ARM_WIDTH 1.0
`define ARM_SETUP_TIME 1.0
`define ARM_HOLD_TIME 0.5
`define ARM_RECOVERY_TIME 1.0
`define ARM_REMOVAL_TIME 0.5

`timescale 1ns/1ps

`ifdef POWER_PINS
`timescale 1ns/1ps
`celldefine
module ADDFH_X1_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(S_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X2_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(S_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X4_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(S_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X8_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(S_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_XL_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(S_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X1_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X2_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X4_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X8_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_XL_A7TULL ( CO, S,VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X1_A7TULL ( CO, S,VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X2_A7TULL ( CO, S,VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X4_A7TULL ( CO, S,VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X8_A7TULL ( CO, S,VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X12_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X2_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X4_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X6_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X8_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X12_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X1_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X2_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X4_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X6_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X8_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_XL_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X12_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X1_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X2_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X4_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X6_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X8_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_XL_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ANTENNA_A7TULL (A,VDD, VSS);
inout VDD, VSS;
input A;

specify

endspecify
endmodule // ANTENNA_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X1_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X2_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X4_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X8_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_XL_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X8_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2B_X1_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1N);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1N;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2B_X2_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1N);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1N;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2B_X4_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1N);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1N;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2B_XL_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1N);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1N;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2_X1_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2_X2_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2_X4_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2_XL_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X1_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X2_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X4_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X8_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_XL_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (out_temp,outA,outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X1_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X2_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X3_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X4_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X6_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X8_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_XL_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_X1_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_X2_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_X4_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_X8_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_XL_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_X1_A7TULL (Y,VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_X2_A7TULL (Y,VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_X4_A7TULL (Y,VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_X8_A7TULL (Y,VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_XL_A7TULL (Y,VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_X1_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_X2_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_X4_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_X8_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_XL_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X1_A7TULL (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X2_A7TULL (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X4_A7TULL (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_XL_A7TULL (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X1_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X2_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X4_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_XL_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33_X1_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33_X2_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33_X4_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33_XL_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X10_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X10_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X12_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X14_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X14_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X16_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X18_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X18_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X20_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X24_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X32_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X4_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X5_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X5_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X6_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X8_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X12_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X16_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X2_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X3_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X4_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X6_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X8_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X12_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X16_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X1_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X20_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X24_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X2_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X32_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X3_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X40_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X40_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X4_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X6_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X8_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X12_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X16_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X1_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X20_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X24_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X2_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X32_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X3_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X40_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X40_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X4_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X6_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X8_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X12_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X16_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X2_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X3_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X4_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X6_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X8_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X12_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X16_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X2_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X4_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X8_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X12_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X16_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X2_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X4_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X8_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DFFHQN_X1_A7TULL (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQN_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQN_X2_A7TULL (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQN_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQN_X4_A7TULL (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQN_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQN_X8_A7TULL (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQN_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQ_X1_A7TULL (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQ_X2_A7TULL (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQ_X4_A7TULL (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQ_X8_A7TULL (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFH_X1_A7TULL (Q, QN,VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFH_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFH_X2_A7TULL (Q, QN,VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFH_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFH_X4_A7TULL (Q, QN,VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFH_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFH_X8_A7TULL (Q, QN,VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFH_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNH_X1_A7TULL (Q, QN,VDD, VSS, CKN, D);
inout VDD, VSS;
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not      IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNH_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNH_X2_A7TULL (Q, QN,VDD, VSS, CKN, D);
inout VDD, VSS;
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not      IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNH_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNH_X4_A7TULL (Q, QN,VDD, VSS, CKN, D);
inout VDD, VSS;
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not      IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNH_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNH_X8_A7TULL (Q, QN,VDD, VSS, CKN, D);
inout VDD, VSS;
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not      IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNH_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRH_X1_A7TULL (Q, QN,VDD, VSS, CKN, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRH_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRH_X2_A7TULL (Q, QN,VDD, VSS, CKN, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRH_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRH_X4_A7TULL (Q, QN,VDD, VSS, CKN, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRH_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRH_X8_A7TULL (Q, QN,VDD, VSS, CKN, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRH_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X1_A7TULL (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X2_A7TULL (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X4_A7TULL (QN,VDD, VSS, CK, D);
inout VDD, VSS;
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X1_A7TULL (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X2_A7TULL (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X4_A7TULL (Q,VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQ_X1_A7TULL (Q,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQ_X2_A7TULL (Q,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQ_X4_A7TULL (Q,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQ_X8_A7TULL (Q,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRQ_X1_A7TULL (Q,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRQ_X2_A7TULL (Q,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRQ_X4_A7TULL (Q,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFR_X1_A7TULL (Q, QN,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFR_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFR_X2_A7TULL (Q, QN,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFR_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFR_X4_A7TULL (Q, QN,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFR_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQ_X1_A7TULL (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQ_X2_A7TULL (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQ_X4_A7TULL (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQ_X8_A7TULL (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X1_A7TULL (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X2_A7TULL (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X4_A7TULL (Q,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQ_X1_A7TULL (Q,VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSRHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQ_X2_A7TULL (Q,VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSRHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQ_X4_A7TULL (Q,VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSRHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQ_X8_A7TULL (Q,VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSRHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSR_X1_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSR_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSR_X2_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSR_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSR_X4_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSR_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFS_X1_A7TULL (Q, QN,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFS_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFS_X2_A7TULL (Q, QN,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFS_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFS_X4_A7TULL (Q, QN,VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFS_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTR_X1_A7TULL (Q, QN,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft_PWR  I0 (n0, dD, clk, dRN, dSN, dEN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTR_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTR_X2_A7TULL (Q, QN,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft_PWR  I0 (n0, dD, clk, dRN, dSN, dEN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTR_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTR_X4_A7TULL (Q, QN,VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft_PWR  I0 (n0, dD, clk, dRN, dSN, dEN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTR_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFF_X1_A7TULL (Q, QN,VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFF_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFF_X2_A7TULL (Q, QN,VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFF_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFF_X4_A7TULL (Q, QN,VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, dD, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFF_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DLY1_X1_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY1_X4_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2_X1_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2_X4_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY3_X1_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY3_X4_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X1_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X4_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module EDFFHQ_X1_A7TULL (Q,VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     B1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFHQ_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFHQ_X2_A7TULL (Q,VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     B1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFHQ_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFHQ_X4_A7TULL (Q,VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     B1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFHQ_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFHQ_X8_A7TULL (Q,VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     B1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFHQ_X8_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTR_X1_A7TULL (Q, QN,VDD, VSS, CK, D, E, RN);
inout VDD, VSS;
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTR_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTR_X2_A7TULL (Q, QN,VDD, VSS, CK, D, E, RN);
inout VDD, VSS;
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTR_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTR_X4_A7TULL (Q, QN,VDD, VSS, CK, D, E, RN);
inout VDD, VSS;
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTR_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFF_X1_A7TULL (Q, QN,VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     B1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not      I1 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFF_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFF_X2_A7TULL (Q, QN,VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     B1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not      I1 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFF_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFF_X4_A7TULL (Q, QN,VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, dD, dCK, dRN, dSN, dE, VDD, VSS, NOTIFIER);
  buf     B1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not      I1 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFF_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ENDCAPTIE19_A7TULL (VDD, VSS);
inout VDD, VSS;

endmodule //ENDCAPTIE19_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL16_A7TULL (VDD, VSS);
inout VDD, VSS;
endmodule //FILL16_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL1_A7TULL (VDD, VSS);
inout VDD, VSS;
endmodule //FILL1_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL2_A7TULL (VDD, VSS);
inout VDD, VSS;
endmodule //FILL2_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL32_A7TULL (VDD, VSS);
inout VDD, VSS;
endmodule //FILL32_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL4_A7TULL (VDD, VSS);
inout VDD, VSS;
endmodule //FILL4_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL64_A7TULL (VDD, VSS);
inout VDD, VSS;
endmodule //FILL64_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL8_A7TULL (VDD, VSS);
inout VDD, VSS;
endmodule //FILL8_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP16_A7TULL (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP32_A7TULL (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP4_A7TULL (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP64_A7TULL (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP64_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP8_A7TULL (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLTIE_A7TULL (VDD, VSS);
inout VDD, VSS;
endmodule //FILLTIE_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module HOLD_X1_A7TULL (Y,VDD, VSS);
inout VDD, VSS;
inout Y;

wire io_wire;

  udp_power(weak0,weak1) I0(Y, io_wire, VDD, VSS);
  udp_power I1(io_wire, Y, VDD, VSS);



specify

endspecify
endmodule // HOLD_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X10_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X10_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X12_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X14_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X14_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X16_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X18_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X18_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X20_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X24_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X32_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X4_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X5_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X5_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X6_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X8_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_XL_A7TULL ( Y,VDD, VSS, A );
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MDFFHQ_X1_A7TULL (Q,VDD, VSS, CK, D0, D1, S0);
inout VDD, VSS;
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff_PWR  I1 (n0, nm, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf      I5 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_S0 ;
wire ENABLE_S0 ;
assign ENABLE_NOT_S0 = (!S0) ? 1'b1:1'b0;
assign ENABLE_S0 = (S0) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK, posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
if (D0==1'b0 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MDFFHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module MDFFHQ_X2_A7TULL (Q,VDD, VSS, CK, D0, D1, S0);
inout VDD, VSS;
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff_PWR  I1 (n0, nm, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf      I5 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_S0 ;
wire ENABLE_S0 ;
assign ENABLE_NOT_S0 = (!S0) ? 1'b1:1'b0;
assign ENABLE_S0 = (S0) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK, posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
if (D0==1'b0 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MDFFHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module MDFFHQ_X4_A7TULL (Q,VDD, VSS, CK, D0, D1, S0);
inout VDD, VSS;
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff_PWR  I1 (n0, nm, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf      I5 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_S0 ;
wire ENABLE_S0 ;
assign ENABLE_NOT_S0 = (!S0) ? 1'b1:1'b0;
assign ENABLE_S0 = (S0) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK, posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
if (D0==1'b0 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MDFFHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module MDFFHQ_X8_A7TULL (Q,VDD, VSS, CK, D0, D1, S0);
inout VDD, VSS;
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff_PWR  I1 (n0, nm, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  buf      I5 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_S0 ;
wire ENABLE_S0 ;
assign ENABLE_NOT_S0 = (!S0) ? 1'b1:1'b0;
assign ENABLE_S0 = (S0) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK, posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
if (D0==1'b0 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MDFFHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module MX2_X12_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X1_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X2_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X3_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X4_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X6_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X8_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_XL_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_X1_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, C, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_X2_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, C, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_X4_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, C, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_X8_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, C, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_XL_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, C, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_X1_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_X2_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_X4_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_X8_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_XL_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_X1_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_X2_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_X4_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_X8_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_XL_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X12_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X1_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X2_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X3_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X4_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X6_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X8_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_XL_A7TULL (Y,VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_X1_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_X2_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_X4_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_X8_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_XL_A7TULL (Y,VDD, VSS, A, B, C, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_X1_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_X2_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_X4_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_X8_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_XL_A7TULL (Y,VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X12_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X1_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X2_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X4_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X8_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_XL_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X12_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X5_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X5_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_XL_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X1_A7TULL (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X2_A7TULL (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X4_A7TULL (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_XL_A7TULL (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X12_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X2_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X3_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X4_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X6_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X8_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_XL_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X1_A7TULL (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X2_A7TULL (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X4_A7TULL (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_XL_A7TULL (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X1_A7TULL (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X2_A7TULL (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X4_A7TULL (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_XL_A7TULL (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X12_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X2_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X4_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X6_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X8_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_XL_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X12_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X1_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X2_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X4_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X8_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_XL_A7TULL (Y,VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X12_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X5_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X5_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_XL_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3B_X1_A7TULL (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3B_X2_A7TULL (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3B_X4_A7TULL (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3B_XL_A7TULL (Y,VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X12_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X2_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X4_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X6_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X8_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_XL_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X1_A7TULL (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X2_A7TULL (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X4_A7TULL (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_XL_A7TULL (Y,VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4B_X1_A7TULL (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4B_X2_A7TULL (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4B_X4_A7TULL (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4B_XL_A7TULL (Y,VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X12_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X1_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X2_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X4_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X6_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X8_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_XL_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X1_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X2_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X4_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X8_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_XL_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X8_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X8_A7TULL (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X1_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X2_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X4_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X8_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_XL_A7TULL (Y,VDD, VSS, A0, A1, B0N);
inout VDD, VSS;
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X1_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X2_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X3_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X4_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X6_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X8_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_XL_A7TULL (Y,VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X1_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X2_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X4_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X8_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_XL_A7TULL (Y,VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B11_X1_A7TULL (Y,VDD, VSS, A0, A1N, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1N, B0, C0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, outA, B0, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B11_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B11_X2_A7TULL (Y,VDD, VSS, A0, A1N, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1N, B0, C0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, outA, B0, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B11_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B11_X4_A7TULL (Y,VDD, VSS, A0, A1N, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1N, B0, C0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, outA, B0, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B11_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B11_XL_A7TULL (Y,VDD, VSS, A0, A1N, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1N, B0, C0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, outA, B0, C0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B11_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_X1_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_X2_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_X4_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_X8_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_XL_A7TULL (Y,VDD, VSS, A0, A1N, B0);
inout VDD, VSS;
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_X1_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_X2_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_X4_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_X8_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_XL_A7TULL (Y,VDD, VSS, A0, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1_X1_A7TULL (Y,VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1_X2_A7TULL (Y,VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1_X4_A7TULL (Y,VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1_XL_A7TULL (Y,VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_X1_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_X2_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_X4_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_X8_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_XL_A7TULL (Y,VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X1_A7TULL (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X2_A7TULL (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X4_A7TULL (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_XL_A7TULL (Y,VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32_X1_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32_X2_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32_X4_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32_XL_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33_X1_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33_X2_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33_X4_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33_XL_A7TULL (Y,VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X12_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X2_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X4_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X6_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X8_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X12_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X1_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X2_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X4_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X6_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X8_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X12_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X1_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X2_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X4_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X6_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X8_A7TULL (Y,VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module SDFFHQN_X1_A7TULL (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQN_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQN_X2_A7TULL (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQN_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQN_X4_A7TULL (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQN_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQN_X8_A7TULL (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQN_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQ_X1_A7TULL (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQ_X2_A7TULL (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQ_X4_A7TULL (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQ_X8_A7TULL (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFH_X1_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFH_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFH_X2_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFH_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFH_X4_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFH_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFH_X8_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFH_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNH_X1_A7TULL (Q, QN,VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNH_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNH_X2_A7TULL (Q, QN,VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNH_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNH_X4_A7TULL (Q, QN,VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNH_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNH_X8_A7TULL (Q, QN,VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNH_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRH_X1_A7TULL (Q, QN,VDD, VSS, CKN, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRH_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRH_X2_A7TULL (Q, QN,VDD, VSS, CKN, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRH_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRH_X4_A7TULL (Q, QN,VDD, VSS, CKN, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRH_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRH_X8_A7TULL (Q, QN,VDD, VSS, CKN, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRH_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X1_A7TULL (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X2_A7TULL (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X4_A7TULL (QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X1_A7TULL (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X2_A7TULL (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X4_A7TULL (Q,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQ_X1_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQ_X2_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQ_X4_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQ_X8_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRQ_X1_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRQ_X2_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRQ_X4_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFR_X1_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFR_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFR_X2_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFR_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFR_X4_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFR_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQ_X1_A7TULL (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQ_X2_A7TULL (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQ_X4_A7TULL (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQ_X8_A7TULL (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X1_A7TULL (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X2_A7TULL (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X4_A7TULL (Q,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQ_X1_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSRHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQ_X2_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSRHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQ_X4_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSRHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQ_X8_A7TULL (Q,VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSRHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSR_X1_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSR_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSR_X2_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSR_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSR_X4_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSR_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFS_X1_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFS_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFS_X2_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFS_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFS_X4_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFS_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTR_X1_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER);
   buf        I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
   not        I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTR_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTR_X2_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER);
   buf        I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
   not        I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTR_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTR_X4_A7TULL (Q, QN,VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER);
   buf        I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
   not        I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTR_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFF_X1_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFF_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFF_X2_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFF_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFF_X4_A7TULL (Q, QN,VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff_PWR  I0 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
  not     I72 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFF_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SEDFFHQ_X1_A7TULL (Q,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER);
   buf       I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQ_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQ_X2_A7TULL (Q,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER);
   buf       I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQ_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQ_X4_A7TULL (Q,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER);
   buf       I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQ_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQ_X8_A7TULL (Q,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER);
   buf       I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQ_X8_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTR_X1_A7TULL (Q, QN,VDD, VSS, CK, D, E, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER);
   buf        I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
   not        I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTR_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTR_X2_A7TULL (Q, QN,VDD, VSS, CK, D, E, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER);
   buf        I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
   not        I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTR_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTR_X4_A7TULL (Q, QN,VDD, VSS, CK, D, E, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER);
   buf        I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
   not        I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTR_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFF_X1_A7TULL (Q, QN,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFF_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFF_X2_A7TULL (Q, QN,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFF_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFF_X4_A7TULL (Q, QN,VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, dD, dCK, dRN, dSI, dSE, dE, VDD, VSS, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFF_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SMDFFHQ_X1_A7TULL (Q,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff_PWR  I1 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_S0_AND_NOT_SE ;
wire ENABLE_S0_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_S0_AND_NOT_SE = (!S0&!SE) ? 1'b1:1'b0;
assign ENABLE_S0_AND_NOT_SE = (S0&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SMDFFHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SMDFFHQ_X2_A7TULL (Q,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff_PWR  I1 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_S0_AND_NOT_SE ;
wire ENABLE_S0_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_S0_AND_NOT_SE = (!S0&!SE) ? 1'b1:1'b0;
assign ENABLE_S0_AND_NOT_SE = (S0&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SMDFFHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SMDFFHQ_X4_A7TULL (Q,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff_PWR  I1 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_S0_AND_NOT_SE ;
wire ENABLE_S0_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_S0_AND_NOT_SE = (!S0&!SE) ? 1'b1:1'b0;
assign ENABLE_S0_AND_NOT_SE = (S0&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SMDFFHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SMDFFHQ_X8_A7TULL (Q,VDD, VSS, CK, D0, D1, S0, SE, SI);
inout VDD, VSS;
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff_PWR  I1 (n0, n1, clk, dRN, dSN, VDD, VSS, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;

wire ENABLE_NOT_S0_AND_NOT_SE ;
wire ENABLE_S0_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_S0_AND_NOT_SE = (!S0&!SE) ? 1'b1:1'b0;
assign ENABLE_S0_AND_NOT_SE = (S0&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SMDFFHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module TBUF_X12_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X16_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X1_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X20_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X24_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X2_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X3_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X4_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X6_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X8_A7TULL ( Y,VDD, VSS, A, OE );
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIEHI_A7TULL (Y,VDD, VSS);
inout VDD, VSS;
output Y;

  buf I0(out_temp, 1'b1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify

endspecify
endmodule // TIEHI_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIELO_A7TULL (Y,VDD, VSS);
inout VDD, VSS;
output Y;

  buf I0(out_temp, 1'b0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify

endspecify
endmodule // TIELO_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X12_A7TULL (ECK,VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, dE, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X16_A7TULL (ECK,VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, dE, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X20_A7TULL (ECK,VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, dE, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X2_A7TULL (ECK,VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, dE, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X3_A7TULL (ECK,VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, dE, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X4_A7TULL (ECK,VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, dE, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X6_A7TULL (ECK,VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, dE, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X8_A7TULL (ECK,VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, dE, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSR_X1_A7TULL (Q, QN,VDD, VSS, D, GN, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dGN);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dGN);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSR_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSR_X2_A7TULL (Q, QN,VDD, VSS, D, GN, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dGN);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dGN);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSR_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSR_X4_A7TULL (Q, QN,VDD, VSS, D, GN, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dGN);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dGN);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSR_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X12_A7TULL (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat_PWR  I1 (n0, n1, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, dCK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X16_A7TULL (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat_PWR  I1 (n0, n1, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, dCK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X20_A7TULL (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat_PWR  I1 (n0, n1, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, dCK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X2_A7TULL (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat_PWR  I1 (n0, n1, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, dCK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X3_A7TULL (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat_PWR  I1 (n0, n1, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, dCK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X4_A7TULL (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat_PWR  I1 (n0, n1, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, dCK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X6_A7TULL (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat_PWR  I1 (n0, n1, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, dCK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X8_A7TULL (ECK,VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat_PWR  I1 (n0, n1, dCK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, dCK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATN_X1_A7TULL (Q, QN,VDD, VSS, D, GN);
inout VDD, VSS;
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN,`ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATN_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATN_X2_A7TULL (Q, QN,VDD, VSS, D, GN);
inout VDD, VSS;
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN,`ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATN_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATN_X4_A7TULL (Q, QN,VDD, VSS, D, GN);
inout VDD, VSS;
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN,`ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATN_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSR_X1_A7TULL (Q, QN,VDD, VSS, D, G, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,dG);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSR_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSR_X2_A7TULL (Q, QN,VDD, VSS, D, G, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,dG);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSR_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSR_X4_A7TULL (Q, QN,VDD, VSS, D, G, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,dG);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSR_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLAT_X1_A7TULL (Q, QN,VDD, VSS, D, G);
inout VDD, VSS;
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,dG);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G,`ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLAT_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLAT_X2_A7TULL (Q, QN,VDD, VSS, D, G);
inout VDD, VSS;
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,dG);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G,`ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLAT_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLAT_X4_A7TULL (Q, QN,VDD, VSS, D, G);
inout VDD, VSS;
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (out_temp, n0);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not      I2 (out__temp, n0);
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0))? out__temp : 1'bx;
not  I3(clk,dG);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G,`ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLAT_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X1_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X2_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X4_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X8_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_XL_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X1_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X2_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X4_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X8_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_XL_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X1_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X2_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X3_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X4_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X8_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_XL_A7TULL (Y,VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X1_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X2_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X4_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X8_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_XL_A7TULL (Y,VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_XL_A7TULL
`endcelldefine
`else

`timescale 1ns/1ps
`celldefine
module ADDFH_X1_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X2_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X4_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_X8_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFH_XL_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFH_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X1_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X2_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X4_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_X8_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDF_XL_A7TULL ( CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDF_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X1_A7TULL ( CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X2_A7TULL ( CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X4_A7TULL ( CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDH_X8_A7TULL ( CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDH_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X12_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X1_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X2_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X4_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X6_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2_X8_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X12_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X1_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X2_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X4_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X6_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_X8_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3_XL_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X12_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X1_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X2_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X4_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X6_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_X8_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4_XL_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ANTENNA_A7TULL (A);
input A;

specify

endspecify
endmodule // ANTENNA_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X1_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X2_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X4_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_X8_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO21_XL_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  or I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO21_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X1_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X2_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X4_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_X8_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO22_XL_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO22_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2B_X1_A7TULL (Y, A0, A1N, B0, B1N);
output Y;
input A0, A1N, B0, B1N;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (Y, outA, outB);


specify
if (B0==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2B_X2_A7TULL (Y, A0, A1N, B0, B1N);
output Y;
input A0, A1N, B0, B1N;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (Y, outA, outB);


specify
if (B0==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2B_X4_A7TULL (Y, A0, A1N, B0, B1N);
output Y;
input A0, A1N, B0, B1N;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (Y, outA, outB);


specify
if (B0==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2B_XL_A7TULL (Y, A0, A1N, B0, B1N);
output Y;
input A0, A1N, B0, B1N;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (Y, outA, outB);


specify
if (B0==1'b0 && B1N==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1N==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2_X1_A7TULL (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2_X2_A7TULL (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2_X4_A7TULL (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AO2B2_XL_A7TULL (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AO2B2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X1_A7TULL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X2_A7TULL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_X4_A7TULL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211_XL_A7TULL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X1_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X2_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X4_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_X8_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21B_XL_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X1_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X2_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X3_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X4_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X6_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_X8_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21_XL_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X1_A7TULL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X2_A7TULL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_X4_A7TULL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221_XL_A7TULL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X1_A7TULL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X2_A7TULL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_X4_A7TULL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222_XL_A7TULL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X1_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X2_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_X4_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22_XL_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_X1_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_X2_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_X4_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_X8_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2B1_XL_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2B1_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_X1_A7TULL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_X2_A7TULL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_X4_A7TULL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_X8_A7TULL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1_XL_A7TULL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_X1_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_X2_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_X4_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_X8_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2_XL_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X1_A7TULL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X2_A7TULL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_X4_A7TULL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31_XL_A7TULL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X1_A7TULL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X2_A7TULL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_X4_A7TULL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32_XL_A7TULL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33_X1_A7TULL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33_X2_A7TULL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33_X4_A7TULL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33_XL_A7TULL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X10_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X10_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X12_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X14_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X14_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X16_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X18_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X18_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X20_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X24_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X2_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X32_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X3_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X4_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X5_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X5_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X6_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUF_X8_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUF_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X12_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X16_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X2_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X3_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X4_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X6_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKAND2_X8_A7TULL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKAND2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X12_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X16_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X1_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X20_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X24_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X2_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X32_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X3_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X40_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X40_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X4_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X6_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUF_X8_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUF_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X12_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X16_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X1_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X20_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X24_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X2_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X32_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X3_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X40_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X40_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X4_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X6_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINV_X8_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINV_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X12_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X16_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X2_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X3_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X4_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X6_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKMX2_X8_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKMX2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X12_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X16_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X2_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X4_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKNAND2_X8_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKNAND2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X12_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X16_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X2_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X4_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKXOR2_X8_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKXOR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DFFHQN_X1_A7TULL (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQN_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQN_X2_A7TULL (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQN_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQN_X4_A7TULL (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQN_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQN_X8_A7TULL (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQN_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQ_X1_A7TULL (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQ_X2_A7TULL (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQ_X4_A7TULL (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQ_X8_A7TULL (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFH_X1_A7TULL (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFH_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFH_X2_A7TULL (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFH_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFH_X4_A7TULL (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFH_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFH_X8_A7TULL (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFH_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNH_X1_A7TULL (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not      IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNH_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNH_X2_A7TULL (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not      IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNH_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNH_X4_A7TULL (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not      IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNH_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNH_X8_A7TULL (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not      IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNH_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRH_X1_A7TULL (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRH_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRH_X2_A7TULL (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRH_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRH_X4_A7TULL (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRH_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRH_X8_A7TULL (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRH_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X1_A7TULL (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X2_A7TULL (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQN_X4_A7TULL (QN, CK, D);
output QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQN_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X1_A7TULL (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X2_A7TULL (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFQ_X4_A7TULL (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQ_X1_A7TULL (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQ_X2_A7TULL (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQ_X4_A7TULL (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQ_X8_A7TULL (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRQ_X1_A7TULL (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRQ_X2_A7TULL (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRQ_X4_A7TULL (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFR_X1_A7TULL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFR_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFR_X2_A7TULL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFR_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFR_X4_A7TULL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFR_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQ_X1_A7TULL (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQ_X2_A7TULL (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQ_X4_A7TULL (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQ_X8_A7TULL (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X1_A7TULL (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X2_A7TULL (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSQ_X4_A7TULL (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQ_X1_A7TULL (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSRHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQ_X2_A7TULL (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSRHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQ_X4_A7TULL (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSRHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQ_X8_A7TULL (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // DFFSRHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSR_X1_A7TULL (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSR_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSR_X2_A7TULL (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSR_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSR_X4_A7TULL (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSR_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFS_X1_A7TULL (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFS_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFS_X2_A7TULL (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFS_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFS_X4_A7TULL (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // DFFS_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTR_X1_A7TULL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft I0 (n0, dD, clk, dRN, dSN, dEN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTR_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTR_X2_A7TULL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft I0 (n0, dD, clk, dRN, dSN, dEN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTR_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTR_X4_A7TULL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft I0 (n0, dD, clk, dRN, dSN, dEN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTR_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFF_X1_A7TULL (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFF_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFF_X2_A7TULL (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFF_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFF_X4_A7TULL (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFF_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DLY1_X1_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY1_X4_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2_X1_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2_X4_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY3_X1_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY3_X4_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X1_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4_X4_A7TULL ( Y, A );
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module EDFFHQ_X1_A7TULL (Q, CK, D, E);
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFHQ_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFHQ_X2_A7TULL (Q, CK, D, E);
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFHQ_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFHQ_X4_A7TULL (Q, CK, D, E);
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFHQ_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFHQ_X8_A7TULL (Q, CK, D, E);
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFHQ_X8_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTR_X1_A7TULL (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTR_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTR_X2_A7TULL (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTR_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTR_X4_A7TULL (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTR_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFF_X1_A7TULL (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFF_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFF_X2_A7TULL (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFF_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFF_X4_A7TULL (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFF_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module ENDCAPTIE19_A7TULL;

endmodule //ENDCAPTIE19_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL16_A7TULL;
endmodule //FILL16_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL1_A7TULL;
endmodule //FILL1_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL2_A7TULL;
endmodule //FILL2_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL32_A7TULL;
endmodule //FILL32_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL4_A7TULL;
endmodule //FILL4_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL64_A7TULL;
endmodule //FILL64_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL8_A7TULL;
endmodule //FILL8_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP16_A7TULL;

specify

endspecify
endmodule // FILLCAP16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP32_A7TULL;

specify

endspecify
endmodule // FILLCAP32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP4_A7TULL;

specify

endspecify
endmodule // FILLCAP4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP64_A7TULL;

specify

endspecify
endmodule // FILLCAP64_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP8_A7TULL;

specify

endspecify
endmodule // FILLCAP8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLTIE_A7TULL;
endmodule //FILLTIE_A7TULL

`endcelldefine
`timescale 1ns/1ps
`celldefine
module HOLD_X1_A7TULL (Y);
inout Y;

wire io_wire;

  buf(weak0,weak1) I0(Y, io_wire);
  buf I1(io_wire, Y);



specify

endspecify
endmodule // HOLD_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X10_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X10_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X12_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X14_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X14_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X16_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X18_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X18_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X1_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X20_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X24_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X2_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X32_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X32_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X3_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X4_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X5_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X5_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X6_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_X8_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INV_XL_A7TULL ( Y, A );
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INV_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MDFFHQ_X1_A7TULL (Q, CK, D0, D1, S0);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff  I1 (n0, nm, clk, dRN, dSN, NOTIFIER);
  buf      I5 (Q, n0);

wire ENABLE_NOT_S0 ;
wire ENABLE_S0 ;
assign ENABLE_NOT_S0 = (!S0) ? 1'b1:1'b0;
assign ENABLE_S0 = (S0) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK, posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
if (D0==1'b0 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MDFFHQ_X1_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module MDFFHQ_X2_A7TULL (Q, CK, D0, D1, S0);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff  I1 (n0, nm, clk, dRN, dSN, NOTIFIER);
  buf      I5 (Q, n0);

wire ENABLE_NOT_S0 ;
wire ENABLE_S0 ;
assign ENABLE_NOT_S0 = (!S0) ? 1'b1:1'b0;
assign ENABLE_S0 = (S0) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK, posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
if (D0==1'b0 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MDFFHQ_X2_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module MDFFHQ_X4_A7TULL (Q, CK, D0, D1, S0);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff  I1 (n0, nm, clk, dRN, dSN, NOTIFIER);
  buf      I5 (Q, n0);

wire ENABLE_NOT_S0 ;
wire ENABLE_S0 ;
assign ENABLE_NOT_S0 = (!S0) ? 1'b1:1'b0;
assign ENABLE_S0 = (S0) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK, posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
if (D0==1'b0 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MDFFHQ_X4_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module MDFFHQ_X8_A7TULL (Q, CK, D0, D1, S0);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff  I1 (n0, nm, clk, dRN, dSN, NOTIFIER);
  buf      I5 (Q, n0);

wire ENABLE_NOT_S0 ;
wire ENABLE_S0 ;
assign ENABLE_NOT_S0 = (!S0) ? 1'b1:1'b0;
assign ENABLE_S0 = (S0) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0 == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0 == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK, posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
if (D0==1'b0 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b0 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MDFFHQ_X8_A7TULL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module MX2_X12_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X1_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X2_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X3_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X4_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X6_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_X8_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2_XL_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_X1_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(Y, A, B, C, C, S0, S1);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_X2_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(Y, A, B, C, C, S0, S1);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_X4_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(Y, A, B, C, C, S0, S1);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_X8_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(Y, A, B, C, C, S0, S1);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX3_XL_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(Y, A, B, C, C, S0, S1);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_X1_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_X2_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_X4_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_X8_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4_XL_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_X1_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_X2_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_X4_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_X8_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2D_XL_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2D_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X12_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X1_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X2_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X3_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X4_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X6_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_X8_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2_XL_A7TULL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_X1_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_X2_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_X4_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_X8_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI3_XL_A7TULL (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b0)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (C==1'b1)
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_X1_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_X2_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_X4_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_X8_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4_XL_A7TULL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X12_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X1_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X2_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X4_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_X8_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2B_XL_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X12_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X1_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X2_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X3_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X4_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X5_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X5_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X6_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_X8_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2_XL_A7TULL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X1_A7TULL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X2_A7TULL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_X4_A7TULL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3B_XL_A7TULL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X12_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X1_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X2_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X3_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X4_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X6_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_X8_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3_XL_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X1_A7TULL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X2_A7TULL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_X4_A7TULL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BB_XL_A7TULL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BB_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X1_A7TULL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X2_A7TULL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_X4_A7TULL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4B_XL_A7TULL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X12_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X1_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X2_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X4_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X6_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_X8_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4_XL_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X12_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X1_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X2_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X4_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_X8_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2B_XL_A7TULL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X12_A7TULL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X1_A7TULL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X2_A7TULL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X3_A7TULL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X4_A7TULL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X5_A7TULL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X5_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X6_A7TULL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_X8_A7TULL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2_XL_A7TULL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3B_X1_A7TULL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3B_X2_A7TULL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3B_X4_A7TULL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3B_XL_A7TULL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X12_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X1_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X2_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X4_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X6_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_X8_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3_XL_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X1_A7TULL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X2_A7TULL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_X4_A7TULL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BB_XL_A7TULL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BB_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4B_X1_A7TULL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4B_X2_A7TULL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4B_X4_A7TULL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4B_XL_A7TULL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X12_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X1_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X2_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X4_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X6_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_X8_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4_XL_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X1_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X2_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X4_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_X8_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA21_XL_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA21_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X1_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X2_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X4_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_X8_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OA22_XL_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OA22_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X1_A7TULL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X2_A7TULL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X4_A7TULL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_X8_A7TULL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211_XL_A7TULL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X1_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X2_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X4_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_X8_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21B_XL_A7TULL (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;



  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21B_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X1_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X2_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X3_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X4_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X6_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_X8_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21_XL_A7TULL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X1_A7TULL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X2_A7TULL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_X4_A7TULL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221_XL_A7TULL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X1_A7TULL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X2_A7TULL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_X4_A7TULL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222_XL_A7TULL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X1_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X2_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X4_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_X8_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22_XL_A7TULL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B11_X1_A7TULL (Y, A0, A1N, B0, C0);
output Y;
input A0, A1N, B0, C0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, outA, B0, C0);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B11_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B11_X2_A7TULL (Y, A0, A1N, B0, C0);
output Y;
input A0, A1N, B0, C0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, outA, B0, C0);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B11_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B11_X4_A7TULL (Y, A0, A1N, B0, C0);
output Y;
input A0, A1N, B0, C0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, outA, B0, C0);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B11_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B11_XL_A7TULL (Y, A0, A1N, B0, C0);
output Y;
input A0, A1N, B0, C0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, outA, B0, C0);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B11_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_X1_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_X2_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_X4_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_X8_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B1_XL_A7TULL (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B1_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_X1_A7TULL (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_X2_A7TULL (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_X4_A7TULL (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_X8_A7TULL (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2B2_XL_A7TULL (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;



  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2B2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1_X1_A7TULL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1_X2_A7TULL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1_X4_A7TULL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1_XL_A7TULL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_X1_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_X2_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_X4_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_X8_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2_XL_A7TULL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X1_A7TULL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X2_A7TULL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_X4_A7TULL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31_XL_A7TULL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32_X1_A7TULL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32_X2_A7TULL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32_X4_A7TULL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32_XL_A7TULL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33_X1_A7TULL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33_X2_A7TULL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33_X4_A7TULL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33_XL_A7TULL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X12_A7TULL (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X1_A7TULL (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X2_A7TULL (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X4_A7TULL (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X6_A7TULL (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2_X8_A7TULL (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X12_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X1_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X2_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X4_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X6_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3_X8_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X12_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X1_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X2_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X4_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X6_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4_X8_A7TULL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module SDFFHQN_X1_A7TULL (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQN_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQN_X2_A7TULL (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQN_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQN_X4_A7TULL (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQN_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQN_X8_A7TULL (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQN_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQ_X1_A7TULL (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQ_X2_A7TULL (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQ_X4_A7TULL (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQ_X8_A7TULL (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFH_X1_A7TULL (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFH_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFH_X2_A7TULL (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFH_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFH_X4_A7TULL (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFH_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFH_X8_A7TULL (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFH_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNH_X1_A7TULL (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNH_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNH_X2_A7TULL (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNH_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNH_X4_A7TULL (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNH_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNH_X8_A7TULL (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNH_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRH_X1_A7TULL (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRH_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRH_X2_A7TULL (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRH_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRH_X4_A7TULL (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRH_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRH_X8_A7TULL (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dD);
$recrem(posedge RN, negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCKN);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSE);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCKN,dSI);
$recrem(posedge SN, negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCKN);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRH_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X1_A7TULL (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X2_A7TULL (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQN_X4_A7TULL (QN, CK, D, SE, SI);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQN_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X1_A7TULL (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X2_A7TULL (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFQ_X4_A7TULL (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQ_X1_A7TULL (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQ_X2_A7TULL (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQ_X4_A7TULL (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQ_X8_A7TULL (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRQ_X1_A7TULL (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRQ_X2_A7TULL (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRQ_X4_A7TULL (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFR_X1_A7TULL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFR_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFR_X2_A7TULL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFR_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFR_X4_A7TULL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFR_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQ_X1_A7TULL (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQ_X2_A7TULL (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQ_X4_A7TULL (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQ_X8_A7TULL (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X1_A7TULL (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X2_A7TULL (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSQ_X4_A7TULL (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQ_X1_A7TULL (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSRHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQ_X2_A7TULL (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSRHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQ_X4_A7TULL (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSRHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQ_X8_A7TULL (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);

endspecify
endmodule // SDFFSRHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSR_X1_A7TULL (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSR_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSR_X2_A7TULL (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSR_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSR_X4_A7TULL (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$recrem(posedge RN, posedge CK &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dCK);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSR_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFS_X1_A7TULL (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFS_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFS_X2_A7TULL (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFS_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFS_X4_A7TULL (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_SE_AND_SN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$recrem(posedge SN, posedge CK, `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dCK);
$width(negedge SN,`ARM_WIDTH,0,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFS_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTR_X1_A7TULL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTR_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTR_X2_A7TULL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTR_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTR_X4_A7TULL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTR_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFF_X1_A7TULL (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFF_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFF_X2_A7TULL (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFF_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFF_X4_A7TULL (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFF_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SEDFFHQ_X1_A7TULL (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQ_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQ_X2_A7TULL (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQ_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQ_X4_A7TULL (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQ_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQ_X8_A7TULL (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQ_X8_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTR_X1_A7TULL (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTR_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTR_X2_A7TULL (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTR_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTR_X4_A7TULL (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dRN);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (0, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, 0);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTR_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFF_X1_A7TULL (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFF_X1_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFF_X2_A7TULL (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFF_X2_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFF_X4_A7TULL (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFF_X4_A7TULL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SMDFFHQ_X1_A7TULL (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff I1 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (Q, n0);

wire ENABLE_NOT_S0_AND_NOT_SE ;
wire ENABLE_S0_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_S0_AND_NOT_SE = (!S0&!SE) ? 1'b1:1'b0;
assign ENABLE_S0_AND_NOT_SE = (S0&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SMDFFHQ_X1_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SMDFFHQ_X2_A7TULL (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff I1 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (Q, n0);

wire ENABLE_NOT_S0_AND_NOT_SE ;
wire ENABLE_S0_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_S0_AND_NOT_SE = (!S0&!SE) ? 1'b1:1'b0;
assign ENABLE_S0_AND_NOT_SE = (S0&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SMDFFHQ_X2_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SMDFFHQ_X4_A7TULL (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff I1 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (Q, n0);

wire ENABLE_NOT_S0_AND_NOT_SE ;
wire ENABLE_S0_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_S0_AND_NOT_SE = (!S0&!SE) ? 1'b1:1'b0;
assign ENABLE_S0_AND_NOT_SE = (S0&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SMDFFHQ_X4_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SMDFFHQ_X8_A7TULL (Q, CK, D0, D1, S0, SE, SI);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff I1 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (Q, n0);

wire ENABLE_NOT_S0_AND_NOT_SE ;
wire ENABLE_S0_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_SE ;
assign ENABLE_NOT_S0_AND_NOT_SE = (!S0&!SE) ? 1'b1:1'b0;
assign ENABLE_S0_AND_NOT_SE = (S0&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,0,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), posedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_NOT_S0_AND_NOT_SE == 1'b1), negedge D0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD0);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), posedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_S0_AND_NOT_SE == 1'b1), negedge D1, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dD1);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge S0, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dS0);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSI);
if (D0==1'b0 && D1==1'b0 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b0 && S0==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b0 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && SE==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b0 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b0 && S0==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b1 || D0==1'b0 && D1==1'b1 && S0==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && D1==1'b1 && S0==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D0==1'b1 && S0==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D1==1'b1 && S0==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SMDFFHQ_X8_A7TULL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module TBUF_X12_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X16_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X1_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X20_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X24_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X24_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X2_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X3_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X4_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X6_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUF_X8_A7TULL ( Y, A, OE );
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (0, 0,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUF_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIEHI_A7TULL (Y);
output Y;

  buf I0(Y, 1'b1);


specify

endspecify
endmodule // TIEHI_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIELO_A7TULL (Y);
output Y;

  buf I0(Y, 1'b0);


specify

endspecify
endmodule // TIELO_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X12_A7TULL (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X16_A7TULL (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X20_A7TULL (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X2_A7TULL (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X3_A7TULL (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X4_A7TULL (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X6_A7TULL (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCA_X8_A7TULL (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);

endspecify
endmodule // TLATNCA_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSR_X1_A7TULL (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dGN);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dGN);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSR_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSR_X2_A7TULL (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dGN);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dGN);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSR_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSR_X4_A7TULL (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dGN);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dGN);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSR_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X12_A7TULL (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X12_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X16_A7TULL (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X16_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X20_A7TULL (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X20_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X2_A7TULL (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X3_A7TULL (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X4_A7TULL (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X6_A7TULL (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X6_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCA_X8_A7TULL (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (0, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dE);
$setuphold(posedge CK, posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);
$setuphold(posedge CK, negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dCK,dSE);

endspecify
endmodule // TLATNTSCA_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATN_X1_A7TULL (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN,`ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATN_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATN_X2_A7TULL (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN,`ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATN_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATN_X4_A7TULL (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dGN,dD);
$width(negedge GN,`ARM_WIDTH,0,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATN_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSR_X1_A7TULL (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,dG);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSR_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSR_X2_A7TULL (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,dG);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSR_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSR_X4_A7TULL (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, dSN);
buf       XX1 (xRN, dRN);

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,dG);

wire ENABLE_RN_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dRN,dG);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER, , ,dSN,dG);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dRN,dSN);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(negedge RN *> (Q +: 1'b0))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, 0);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b1 && G==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, 0);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(negedge SN *> (QN -: 1'b1))=(0, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSR_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLAT_X1_A7TULL (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,dG);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G,`ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLAT_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLAT_X2_A7TULL (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,dG);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G,`ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLAT_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLAT_X4_A7TULL (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,dG);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER, , ,dG,dD);
$width(posedge G,`ARM_WIDTH,0,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLAT_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X1_A7TULL (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X2_A7TULL (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X4_A7TULL (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_X8_A7TULL (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2_XL_A7TULL (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X1_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X2_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X4_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_X8_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3_XL_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X1_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X2_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X3_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X3_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X4_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_X8_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2_XL_A7TULL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2_XL_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X1_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X1_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X2_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X2_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X4_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X4_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_X8_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_X8_A7TULL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3_XL_A7TULL (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3_XL_A7TULL
`endcelldefine
`endif
