library verilog;
use verilog.vl_types.all;
entity aftab_DARU_TB is
end aftab_DARU_TB;
